
module problem_9_11(
    input [7:0] data_in,
    output [7:0] data_out,
    input push,
    input pop,
    input clk,
    input reset,
    output full,
    output empty
    );


endmodule
