-- ==========================
-- Listing 2.1 Even detector
-- ==========================

library ieee;
use ieee.std_logic_1164.all;

-- entity declaration
entity even_detector is
	port(
		a: in std_logic_vector(2 downto 0);
		b: in std_logic_vector(2 downto 0);
		even: out std_logic;
		odd:	out std_logic
	);
end even_detector;

-- architecture body
architecture sop_arch of even_detector is
	signal p1, p2, p3, p4, q1, q2, q3, q4 : std_logic;
begin
	even 	<= (p1 or p2) or (p3 or p4) 						after 20 ns;
	p1		<= (not a(2)) and (not a(1)) and (not a(0)) 	after 15 ns;
	p2		<= (not a(2)) and a(1) and a(0) 					after 12 ns;
	p3		<= a(2) and (not a(1)) and a(0)					after 12 ns;
	p4		<= a(2) and a(1) and (not a(0))					after 12 ns;

	odd 	<= not ((q1 or q2) or (q3 or q4))				after 20 ns;
	q1		<= (not b(2)) and (not b(1)) and (not b(0)) 	after 15 ns;
	q2		<= (not b(2)) and b(1) and b(0) 					after 12 ns;
	q3		<= b(2) and (not b(1)) and b(0)					after 12 ns;
	q4		<= b(2) and b(1) and (not b(0))					after 12 ns;
end sop_arch;